/*
Create a class "my_object" by extending the UVM_OBJECT class. Add three logic datatype datamembers "a", "b", and "c" with sizes of 2, 4, and 8 respectively. Generate a random value for all the data members and send the values of the variables to the console by using the print method.
*/

class className extends superClass;
  function new();
    
  endfunction //new()
endclass //className extends superClass